library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bcd_decoder is
  port (
	 bcd_num       : in  std_logic_vector(31 downto 0);
    seven_seg_num : out std_logic_vector(31 downto 0)
  );
end entity;

architecture arch of bcd_decoder is
begin
  process ( bcd_num ) begin
	case bcd_num is
   when "00000000000000000000000000000000" => seven_seg_num <= not ("1111110" & "1111110" & "000000000000000000"); -- 00
   when "00000000000000000000000000000001" => seven_seg_num <= not ("1111110" & "0000110" & "000000000000000000"); -- 01
   when "00000000000000000000000000000010" => seven_seg_num <= not ("1111110" & "1101101" & "000000000000000000"); -- 02
   when "00000000000000000000000000000011" => seven_seg_num <= not ("1111110" & "1111001" & "000000000000000000"); -- 03
   when "00000000000000000000000000000100" => seven_seg_num <= not ("1111110" & "0110011" & "000000000000000000"); -- 04
   when "00000000000000000000000000000101" => seven_seg_num <= not ("1111110" & "1011011" & "000000000000000000"); -- 05
   when "00000000000000000000000000000110" => seven_seg_num <= not ("1111110" & "1011111" & "000000000000000000"); -- 06
   when "00000000000000000000000000000111" => seven_seg_num <= not ("1111110" & "1110000" & "000000000000000000"); -- 07
   when "00000000000000000000000000001000" => seven_seg_num <= not ("1111110" & "1111111" & "000000000000000000"); -- 08
   when "00000000000000000000000000001001" => seven_seg_num <= not ("1111110" & "1111011" & "000000000000000000"); -- 09

   when "00000000000000000000000000001010" => seven_seg_num <= not ("0000110" & "1111110" & "000000000000000000"); -- 10
   when "00000000000000000000000000001011" => seven_seg_num <= not ("0000110" & "0000110" & "000000000000000000"); -- 11
   when "00000000000000000000000000001100" => seven_seg_num <= not ("0000110" & "1101101" & "000000000000000000"); -- 12
   when "00000000000000000000000000001101" => seven_seg_num <= not ("0000110" & "1111001" & "000000000000000000"); -- 13
   when "00000000000000000000000000001110" => seven_seg_num <= not ("0000110" & "0110011" & "000000000000000000"); -- 14
   when "00000000000000000000000000001111" => seven_seg_num <= not ("0000110" & "1011011" & "000000000000000000"); -- 15
   when "00000000000000000000000000010000" => seven_seg_num <= not ("0000110" & "1011111" & "000000000000000000"); -- 16
   when "00000000000000000000000000010001" => seven_seg_num <= not ("0000110" & "1110000" & "000000000000000000"); -- 17
   when "00000000000000000000000000010010" => seven_seg_num <= not ("0000110" & "1111111" & "000000000000000000"); -- 18
   when "00000000000000000000000000010011" => seven_seg_num <= not ("0000110" & "1111011" & "000000000000000000"); -- 19

   when "00000000000000000000000000010100" => seven_seg_num <= not ("1101101" & "1111110" & "000000000000000000"); -- 20
   when "00000000000000000000000000010101" => seven_seg_num <= not ("1101101" & "0000110" & "000000000000000000"); -- 21
   when "00000000000000000000000000010110" => seven_seg_num <= not ("1101101" & "1101101" & "000000000000000000"); -- 22
   when "00000000000000000000000000010111" => seven_seg_num <= not ("1101101" & "1111001" & "000000000000000000"); -- 23
   when "00000000000000000000000000011000" => seven_seg_num <= not ("1101101" & "0110011" & "000000000000000000"); -- 24
   when "00000000000000000000000000011001" => seven_seg_num <= not ("1101101" & "1011011" & "000000000000000000"); -- 25
   when "00000000000000000000000000011010" => seven_seg_num <= not ("1101101" & "1011111" & "000000000000000000"); -- 26
   when "00000000000000000000000000011011" => seven_seg_num <= not ("1101101" & "1110000" & "000000000000000000"); -- 27
   when "00000000000000000000000000011100" => seven_seg_num <= not ("1101101" & "1111111" & "000000000000000000"); -- 28
   when "00000000000000000000000000011101" => seven_seg_num <= not ("1101101" & "1111011" & "000000000000000000"); -- 29

   when "00000000000000000000000000011110" => seven_seg_num <= not ("1111001" & "1111110" & "000000000000000000"); -- 30
   when "00000000000000000000000000011111" => seven_seg_num <= not ("1111001" & "0000110" & "000000000000000000"); -- 31
   when "00000000000000000000000000100000" => seven_seg_num <= not ("1111001" & "1101101" & "000000000000000000"); -- 32
   when "00000000000000000000000000100001" => seven_seg_num <= not ("1111001" & "1111001" & "000000000000000000"); -- 33
   when "00000000000000000000000000100010" => seven_seg_num <= not ("1111001" & "0110011" & "000000000000000000"); -- 34
   when "00000000000000000000000000100011" => seven_seg_num <= not ("1111001" & "1011011" & "000000000000000000"); -- 35
   when "00000000000000000000000000100100" => seven_seg_num <= not ("1111001" & "1011111" & "000000000000000000"); -- 36
   when "00000000000000000000000000100101" => seven_seg_num <= not ("1111001" & "1110000" & "000000000000000000"); -- 37
   when "00000000000000000000000000100110" => seven_seg_num <= not ("1111001" & "1111111" & "000000000000000000"); -- 38
   when "00000000000000000000000000100111" => seven_seg_num <= not ("1111001" & "1111011" & "000000000000000000"); -- 39

   when "00000000000000000000000000101000" => seven_seg_num <= not ("0110011" & "1111110" & "000000000000000000"); -- 40
   when "00000000000000000000000000101001" => seven_seg_num <= not ("0110011" & "0000110" & "000000000000000000"); -- 41
   when "00000000000000000000000000101010" => seven_seg_num <= not ("0110011" & "1101101" & "000000000000000000"); -- 42
   when "00000000000000000000000000101011" => seven_seg_num <= not ("0110011" & "1111001" & "000000000000000000"); -- 43
   when "00000000000000000000000000101100" => seven_seg_num <= not ("0110011" & "0110011" & "000000000000000000"); -- 44
   when "00000000000000000000000000101101" => seven_seg_num <= not ("0110011" & "1011011" & "000000000000000000"); -- 45
   when "00000000000000000000000000101110" => seven_seg_num <= not ("0110011" & "1011111" & "000000000000000000"); -- 46
   when "00000000000000000000000000101111" => seven_seg_num <= not ("0110011" & "1110000" & "000000000000000000"); -- 47
   when "00000000000000000000000000110000" => seven_seg_num <= not ("0110011" & "1111111" & "000000000000000000"); -- 48
   when "00000000000000000000000000110001" => seven_seg_num <= not ("0110011" & "1111011" & "000000000000000000"); -- 49

   when "00000000000000000000000000110010" => seven_seg_num <= not ("1011011" & "1111110" & "000000000000000000"); -- 50
   when "00000000000000000000000000110011" => seven_seg_num <= not ("1011011" & "0000110" & "000000000000000000"); -- 51
   when "00000000000000000000000000110100" => seven_seg_num <= not ("1011011" & "1101101" & "000000000000000000"); -- 52
   when "00000000000000000000000000110101" => seven_seg_num <= not ("1011011" & "1111001" & "000000000000000000"); -- 53
   when "00000000000000000000000000110110" => seven_seg_num <= not ("1011011" & "0110011" & "000000000000000000"); -- 54
   when "00000000000000000000000000110111" => seven_seg_num <= not ("1011011" & "1011011" & "000000000000000000"); -- 55
   when "00000000000000000000000000111000" => seven_seg_num <= not ("1011011" & "1011111" & "000000000000000000"); -- 56
   when "00000000000000000000000000111001" => seven_seg_num <= not ("1011011" & "1110000" & "000000000000000000"); -- 57
   when "00000000000000000000000000111010" => seven_seg_num <= not ("1011011" & "1111111" & "000000000000000000"); -- 58
   when "00000000000000000000000000111011" => seven_seg_num <= not ("1011011" & "1111011" & "000000000000000000"); -- 59
   when others                             => seven_seg_num <= not ("1011110" & "1011110" & "000000000000000000"); --  Else muestre GG
  end case;
  end process;
end architecture;
